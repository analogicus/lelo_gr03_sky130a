*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/BANDGAP_CIRCUIT_TB_lpe.spi
#else
.include ../../../work/xsch/BANDGAP_CIRCUIT_TB.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
VPTAT I_PTAT VSS 0.5

.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0

*ptran 0 0 0 1n 1u 0

#ifdef Nosweep
tran 10n {t_stop}
write {cicname}.raw
#else
set fend = .raw
foreach vtemp {temperatures}
  option temp=$vtemp
  tran 10n {t_stop}
  write {cicname}_$vtemp$fend
end

#endif

quit


.endc

.end