*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/BANDGAP_OTA_lpe.spi
#else
.include ../../../work/xsch/BANDGAP_OTA.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}    

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
* VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VDD VDD_1V8 VSS dc {AVDD}

*INPUT SIGNALS
VPWR_ON PWR_ON VSS dc 0

VINP INP VSS SIN(0.6 5m 1Meg)
VINN INN VSS SIN(0.6 -5m 1Meg)


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

* --- Operating point ---
op
save all
write op.raw

* --- ________________ ---

optran 0 0 0 1n 1u 0


tran 1n 5u 1p
write
quit


.endc

.end
