** sch_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/LELO_GR03_SKY130A/BANDGAP_OTA_TB.sch
**.subckt BANDGAP_OTA_TB
xdut net2 net3 net3 net1 0 BANDGAP_OTA
xcap net1 0 JNWTR_CAPX1
V1 net2 0 1.8
V2 net3 0 0.6
**** begin user architecture code


.param mc_mm_switch=0
.param mc_pr_switch=0

.lib ../../../tech/ngspice/temperature.spi Tl
.lib ../../../tech/ngspice/corners.spi Kss
.lib ../../../tech/ngspice/supply.spi Vl
.include ../../../../cpdk/ngspice/ideal_circuits.spi

.option SEED=1
.option savecurrents
.control
set interactive
optran 0 0 0 10n 1u 0
save all
save @m.xdut.*.xm1.msky130_fd_pr__*[id]
save @m.xdut.*.xm1.msky130_fd_pr__*[gm]
save @m.xdut.*.xm1.msky130_fd_pr__*[vth]
save @m.xdut.*.xm1.msky130_fd_pr__*[vdsat]
op
write BANDGAP_OTA_TB.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  LELO_GR03_SKY130A/BANDGAP_OTA.sym # of pins=5
** sym_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/LELO_GR03_SKY130A/BANDGAP_OTA.sym
** sch_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/LELO_GR03_SKY130A/BANDGAP_OTA.sch
.subckt BANDGAP_OTA VDD IN- IN+ OUT VSS
*.ipin VDD
*.ipin VSS
*.opin OUT
*.ipin IN+
*.ipin IN-
x8<4> net2<4> net1 VDD VDD JNWATR_PCH_4C5F0
x8<3> net2<3> net1 VDD VDD JNWATR_PCH_4C5F0
x8<2> net2<2> net1 VDD VDD JNWATR_PCH_4C5F0
x8<1> net2<1> net1 VDD VDD JNWATR_PCH_4C5F0
x8<0> net2<0> net1 VDD VDD JNWATR_PCH_4C5F0
x2 net1 net1 VDD VDD JNWATR_PCH_4C5F0
x3 net1 net4 VSS JNWTR_RPPO16
x2<4> OUT IN- net2<4> VDD JNWATR_PCH_4C5F0
x2<3> OUT IN- net2<3> VDD JNWATR_PCH_4C5F0
x2<2> OUT IN- net2<2> VDD JNWATR_PCH_4C5F0
x2<1> OUT IN- net2<1> VDD JNWATR_PCH_4C5F0
x2<0> OUT IN- net2<0> VDD JNWATR_PCH_4C5F0
x3<4> net3 IN+ net2<4> VDD JNWATR_PCH_4C5F0
x3<3> net3 IN+ net2<3> VDD JNWATR_PCH_4C5F0
x3<2> net3 IN+ net2<2> VDD JNWATR_PCH_4C5F0
x3<1> net3 IN+ net2<1> VDD JNWATR_PCH_4C5F0
x3<0> net3 IN+ net2<0> VDD JNWATR_PCH_4C5F0
x6 net4 VSS VSS JNWTR_RPPO16
x1 net5 net3 VSS VSS JNWATR_NCH_4C5F0
x4 net6 net3 VSS VSS JNWATR_NCH_4C5F0
x5 net3 net3 net6 VSS JNWATR_NCH_4C5F0
x7 OUT net3 net5 VSS JNWATR_NCH_4C5F0
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO16.sym # of pins=3
** sym_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sym
** sch_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sch
.subckt JNWTR_RPPO16 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES16
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES16.sym # of pins=3
** sym_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sym
** sch_path: /home/kim/pro/aicex/ip/lelo_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sch
.subckt JNWTR_RES16 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 INT_7 INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_8 INT_8 INT_7 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_9 INT_9 INT_8 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_10 INT_10 INT_9 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_11 INT_11 INT_10 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_12 INT_12 INT_11 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_13 INT_13 INT_12 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_14 INT_14 INT_13 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_15 P INT_14 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
